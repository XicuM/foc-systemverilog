`timescale 1ns / 1ps

module inverter #(
    
)(
    input logic clk, en, nrst,
    input logic [] gates,
    output logic [] v_phases
);

endmodule